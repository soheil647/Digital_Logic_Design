library verilog;
use verilog.vl_types.all;
entity TB_Sin is
end TB_Sin;
