library verilog;
use verilog.vl_types.all;
entity testQ is
end testQ;
